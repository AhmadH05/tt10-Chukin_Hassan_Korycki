/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */


`default_nettype none

module tt_um_my_adder (  
    input  wire [7:0] ui_in,    
    output wire [7:0] uo_out,   
    input  wire [7:0] uio_in,   
    output wire [7:0] uio_out,  
    output wire [7:0] uio_oe,   
    input  wire       ena,      
    input  wire       clk,      
    input  wire       rst_n     
);

  assign uo_out = ui_in[3:0] + ui_in[7:4];  

  assign uio_out = 8'b00000000;
  assign uio_oe  = 8'b00000000;

  wire _unused = &{ena, clk, rst_n};

endmodule
